module valve

pub struct ICvar {}
